/*
 * @Author: German Cano Quiveu, germancq@gmail.com 
 * @Date: 2019-09-21 22:20:24 
 * @Last Modified by: German Cano Quiveu, germancq@gmail.com
 * @Last Modified time: 2019-09-21 22:20:56
 */
